module beat32 (
    input wire clk,
    input wire rst,
    output reg count_en
);

wire [4:0] load = 5'b11111;

reg [4:0] next_val;
wire [4:0] val; 
dffr #(.WIDTH(5)) current_val(
.clk (clk), .r (rst), .d (next_val), .q (val)
);

always @(*) begin
    
    case (rst)
        1'b1: begin
            next_val = 0;
        end 
        1'b0: begin
            if (next_val == 5'b0) begin
                count_en = 1'b1;
                next_val = load ;
            end 
            else begin
                count_en = 1'b0;
                next_val = val - 1'b1 ;

            end
       end
     endcase

end
endmodule
